module tb;
	logic [31:0] out [784];
	test test_mod(.weight_data(out));
endmodule