module tb;
	logic out [10];
	Network net(.guess(out));
endmodule