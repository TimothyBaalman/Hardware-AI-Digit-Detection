module tb;
	logic [31:0] out [784];
	test test_mod(.px_data(out));
endmodule