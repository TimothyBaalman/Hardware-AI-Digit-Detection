module multiplier_2c_4b(
	input [3:0] x,
	input [3:0] y,
	output [3:0] result //Shift output by chopping first 2 and last 2 bits.
);
	wire [7:0] output;

	
endmodule