module tb;
	logic [31:0] out;
	Network net(.guess(out));
endmodule