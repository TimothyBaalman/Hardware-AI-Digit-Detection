module tb;
	logic [31:0] out [10];
	Network net(.guess(out));
endmodule