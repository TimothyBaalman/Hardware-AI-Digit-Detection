module tb;
	test test_mod();
endmodule